--*****************************************************************************
--***************************  VHDL Source Code  ******************************
--*****************************************************************************
--
--  DESIGNER NAME:  Andrew Serra
--
--       LAB NAME:  Lab 1 - Introduction
--
--      FILE NAME:  template.vhd
--
-------------------------------------------------------------------------------
--
--  DESCRIPTION
--
--    This design will create a circuit that has a switch  
--    and a LED. If the signal from the switch is high, the 
--    LED will output high. if the switch is low, the LED will
--    be outputting low.
--
-------------------------------------------------------------------------------
--
--  REVISION HISTORY
--
--  _______________________________________________________________________
-- |  DATE    | USER | Ver |  Description                                  |
-- |==========+======+=====+================================================
-- |          |      |     |
-- | 08/29/20 | ACS  | 1.0 | Created
-- |          |      |     |
--
--*****************************************************************************
--*****************************************************************************

------------------------------------------------------------------------------
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
-- ||||                                                                   ||||
-- ||||                    COMPONENT PACKAGE                              ||||
-- ||||                                                                   ||||
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE template_pkg IS
  COMPONENT template IS 
    PORT (
      switch   : IN  std_logic;
      led      : OUT std_logic
      );
  END COMPONENT;
END PACKAGE template_pkg;



------------------------------------------------------------------------------
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
-- |||| 
-- |||| COMPONENT DESCRIPTION 
-- |||| 
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY template IS
  PORT (
      switch   : IN  std_logic;
      led      : OUT  std_logic
    );
END ENTITY template;

ARCHITECTURE behave OF template IS

BEGIN

    led <= '1' WHEN (switch = '1') ELSE '0';

END ARCHITECTURE behave;
