--*****************************************************************************
--***************************  VHDL Source Code  ******************************
--*****************************************************************************
--
--  DESIGNER NAME:  Andrew Serra
--
--       LAB NAME:  Homework 2
--
--      FILE NAME:  and_4.vhd
--
-------------------------------------------------------------------------------
--
--  DESCRIPTION
--
--    This design will produce an AND gate for four inputs. 
--
--
-------------------------------------------------------------------------------
--
--  REVISION HISTORY
--
--  _______________________________________________________________________
-- |  DATE    | USER | Ver |  Description                                  |
-- |==========+======+=====+================================================
-- |          |      |     |
-- | 09/03/20 | ACS  | 1.0 | Created
-- |          |      |     |
--
--*****************************************************************************
--*****************************************************************************

------------------------------------------------------------------------------
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
-- ||||                                                                   ||||
-- ||||                    COMPONENT PACKAGE                              ||||
-- ||||                                                                   ||||
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;

PACKAGE and_4_pkg IS
    COMPONENT and_4 IS
	    PORT (
	        inputs : IN std_logic_vector(3 DOWNTO 0);
		    output : OUT std_logic
	    );
	END COMPONENT;
END PACKAGE and_4_pkg;

------------------------------------------------------------------------------
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
-- |||| 
-- |||| COMPONENT DESCRIPTION 
-- |||| 
-- |||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||||
------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY and_4 IS
    PORT (
		inputs    : IN std_logic_vector(3 DOWNTO 0);
		output    : OUT std_logic
	);
END ENTITY and_4;

ARCHITECTURE behavior OF and_4 IS

BEGIN

    output <= '1' WHEN inputs = "1111" ELSE '0';

END ARCHITECTURE behavior;